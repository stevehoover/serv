../../prepared.sv